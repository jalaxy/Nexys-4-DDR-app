module RegFile(clk, rst, rsc, rtc, rdc, rs, rt, rd, rtin);
    input clk, rst;
    input [4:0] rsc, rtc, rdc;
    output [31:0] rs;
    inout [31:0] rt;
    input [31:0] rd;
    input rtin;

    wire [31:0] ena;
    assign ena = ({31'b0, rtin} << rtc) | (32'b1 << rdc);
    wire [31:0] din[0:31];
    wire [31:0] dout[0:31];
    assign din[0]  = rtc == 5'd0  && rtin ? rt : (rdc == 5'd0  ? rd : 32'bz);
    assign din[1]  = rtc == 5'd1  && rtin ? rt : (rdc == 5'd1  ? rd : 32'bz);
    assign din[2]  = rtc == 5'd2  && rtin ? rt : (rdc == 5'd2  ? rd : 32'bz);
    assign din[3]  = rtc == 5'd3  && rtin ? rt : (rdc == 5'd3  ? rd : 32'bz);
    assign din[4]  = rtc == 5'd4  && rtin ? rt : (rdc == 5'd4  ? rd : 32'bz);
    assign din[5]  = rtc == 5'd5  && rtin ? rt : (rdc == 5'd5  ? rd : 32'bz);
    assign din[6]  = rtc == 5'd6  && rtin ? rt : (rdc == 5'd6  ? rd : 32'bz);
    assign din[7]  = rtc == 5'd7  && rtin ? rt : (rdc == 5'd7  ? rd : 32'bz);
    assign din[8]  = rtc == 5'd8  && rtin ? rt : (rdc == 5'd8  ? rd : 32'bz);
    assign din[9]  = rtc == 5'd9  && rtin ? rt : (rdc == 5'd9  ? rd : 32'bz);
    assign din[10] = rtc == 5'd10 && rtin ? rt : (rdc == 5'd10 ? rd : 32'bz);
    assign din[11] = rtc == 5'd11 && rtin ? rt : (rdc == 5'd11 ? rd : 32'bz);
    assign din[12] = rtc == 5'd12 && rtin ? rt : (rdc == 5'd12 ? rd : 32'bz);
    assign din[13] = rtc == 5'd13 && rtin ? rt : (rdc == 5'd13 ? rd : 32'bz);
    assign din[14] = rtc == 5'd14 && rtin ? rt : (rdc == 5'd14 ? rd : 32'bz);
    assign din[15] = rtc == 5'd15 && rtin ? rt : (rdc == 5'd15 ? rd : 32'bz);
    assign din[16] = rtc == 5'd16 && rtin ? rt : (rdc == 5'd16 ? rd : 32'bz);
    assign din[17] = rtc == 5'd17 && rtin ? rt : (rdc == 5'd17 ? rd : 32'bz);
    assign din[18] = rtc == 5'd18 && rtin ? rt : (rdc == 5'd18 ? rd : 32'bz);
    assign din[19] = rtc == 5'd19 && rtin ? rt : (rdc == 5'd19 ? rd : 32'bz);
    assign din[20] = rtc == 5'd20 && rtin ? rt : (rdc == 5'd20 ? rd : 32'bz);
    assign din[21] = rtc == 5'd21 && rtin ? rt : (rdc == 5'd21 ? rd : 32'bz);
    assign din[22] = rtc == 5'd22 && rtin ? rt : (rdc == 5'd22 ? rd : 32'bz);
    assign din[23] = rtc == 5'd23 && rtin ? rt : (rdc == 5'd23 ? rd : 32'bz);
    assign din[24] = rtc == 5'd24 && rtin ? rt : (rdc == 5'd24 ? rd : 32'bz);
    assign din[25] = rtc == 5'd25 && rtin ? rt : (rdc == 5'd25 ? rd : 32'bz);
    assign din[26] = rtc == 5'd26 && rtin ? rt : (rdc == 5'd26 ? rd : 32'bz);
    assign din[27] = rtc == 5'd27 && rtin ? rt : (rdc == 5'd27 ? rd : 32'bz);
    assign din[28] = rtc == 5'd28 && rtin ? rt : (rdc == 5'd28 ? rd : 32'bz);
    assign din[29] = rtc == 5'd29 && rtin ? rt : (rdc == 5'd29 ? rd : 32'bz);
    assign din[30] = rtc == 5'd30 && rtin ? rt : (rdc == 5'd30 ? rd : 32'bz);
    assign din[31] = rtc == 5'd31 && rtin ? rt : (rdc == 5'd31 ? rd : 32'bz);
    Reg32 r0 (clk, 1,   ena[5'd0],  din[0],  dout[0]);
    Reg32 r1 (clk, rst, ena[5'd1],  din[1],  dout[1]);
    Reg32 r2 (clk, rst, ena[5'd2],  din[2],  dout[2]);
    Reg32 r3 (clk, rst, ena[5'd3],  din[3],  dout[3]);
    Reg32 r4 (clk, rst, ena[5'd4],  din[4],  dout[4]);
    Reg32 r5 (clk, rst, ena[5'd5],  din[5],  dout[5]);
    Reg32 r6 (clk, rst, ena[5'd6],  din[6],  dout[6]);
    Reg32 r7 (clk, rst, ena[5'd7],  din[7],  dout[7]);
    Reg32 r8 (clk, rst, ena[5'd8],  din[8],  dout[8]);
    Reg32 r9 (clk, rst, ena[5'd9],  din[9],  dout[9]);
    Reg32 r10(clk, rst, ena[5'd10], din[10], dout[10]);
    Reg32 r11(clk, rst, ena[5'd11], din[11], dout[11]);
    Reg32 r12(clk, rst, ena[5'd12], din[12], dout[12]);
    Reg32 r13(clk, rst, ena[5'd13], din[13], dout[13]);
    Reg32 r14(clk, rst, ena[5'd14], din[14], dout[14]);
    Reg32 r15(clk, rst, ena[5'd15], din[15], dout[15]);
    Reg32 r16(clk, rst, ena[5'd16], din[16], dout[16]);
    Reg32 r17(clk, rst, ena[5'd17], din[17], dout[17]);
    Reg32 r18(clk, rst, ena[5'd18], din[18], dout[18]);
    Reg32 r19(clk, rst, ena[5'd19], din[19], dout[19]);
    Reg32 r20(clk, rst, ena[5'd20], din[20], dout[20]);
    Reg32 r21(clk, rst, ena[5'd21], din[21], dout[21]);
    Reg32 r22(clk, rst, ena[5'd22], din[22], dout[22]);
    Reg32 r23(clk, rst, ena[5'd23], din[23], dout[23]);
    Reg32 r24(clk, rst, ena[5'd24], din[24], dout[24]);
    Reg32 r25(clk, rst, ena[5'd25], din[25], dout[25]);
    Reg32 r26(clk, rst, ena[5'd26], din[26], dout[26]);
    Reg32 r27(clk, rst, ena[5'd27], din[27], dout[27]);
    Reg32 r28(clk, rst, ena[5'd28], din[28], dout[28]);
    Reg32 r29(clk, rst, ena[5'd29], din[29], dout[29]);
    Reg32 r30(clk, rst, ena[5'd30], din[30], dout[30]);
    Reg32 r31(clk, rst, ena[5'd31], din[31], dout[31]);
    assign rs = dout[rsc];
    assign rt = rtin ? 32'dz : dout[rtc];


    wire [31:0] array_reg[0:31];
    assign array_reg[0]  = dout[5'd0];
    assign array_reg[1]  = dout[5'd1];
    assign array_reg[2]  = dout[5'd2];
    assign array_reg[3]  = dout[5'd3];
    assign array_reg[4]  = dout[5'd4];
    assign array_reg[5]  = dout[5'd5];
    assign array_reg[6]  = dout[5'd6];
    assign array_reg[7]  = dout[5'd7];
    assign array_reg[8]  = dout[5'd8];
    assign array_reg[9]  = dout[5'd9];
    assign array_reg[10] = dout[5'd10];
    assign array_reg[11] = dout[5'd11];
    assign array_reg[12] = dout[5'd12];
    assign array_reg[13] = dout[5'd13];
    assign array_reg[14] = dout[5'd14];
    assign array_reg[15] = dout[5'd15];
    assign array_reg[16] = dout[5'd16];
    assign array_reg[17] = dout[5'd17];
    assign array_reg[18] = dout[5'd18];
    assign array_reg[19] = dout[5'd19];
    assign array_reg[20] = dout[5'd20];
    assign array_reg[21] = dout[5'd21];
    assign array_reg[22] = dout[5'd22];
    assign array_reg[23] = dout[5'd23];
    assign array_reg[24] = dout[5'd24];
    assign array_reg[25] = dout[5'd25];
    assign array_reg[26] = dout[5'd26];
    assign array_reg[27] = dout[5'd27];
    assign array_reg[28] = dout[5'd28];
    assign array_reg[29] = dout[5'd29];
    assign array_reg[30] = dout[5'd30];
    assign array_reg[31] = dout[5'd31];
endmodule

module Reg32(clk, rst, ena, din, dout);
    input clk, rst, ena;
    input [31:0] din;
    output [31:0] dout;

    reg [31:0] data;
    wire clk_ena;
    assign clk_ena = clk & ena;
    assign dout = data;
    always @(posedge clk_ena or posedge rst)
        data = rst ? 32'd0 : din;
endmodule