`define logN 3
`define N 4096
`define M 16
